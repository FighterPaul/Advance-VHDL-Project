

library ieee;
use ieee.std_logic_1164.all;


entity InterfaceLCD is 
port
(
    clk : in std_logic;

    byte_in : in std_logic_vector(127 downto 0);

    lcd_rw : out std_logic;
    lcd_rs : out std_logic;
    lcd_e : out std_logic;
    data_out : out std_logic_vector(7 downto 0)
);
end entity;


architecture arch of InterfaceLCD is

    type arr_command is array(1 to 6) of std_logic_vector(7 downto 0);
    constant command_rom : arr_command := (X"38", X"0C", X"06", X"01", X"C0", X"C0");



    type arr_char is array(1 to 16) of std_logic_vector(7 downto 0);
    constant byte_rom : arr_char := (X"30"X"31"X"32"X"33"X"34"X"35"X"36"X"37", X"38", X"39",
                    X"41"X"42"X"20"X"20"X"20"X"20");

    
    signal en_timing : integer range 0 to 100000 := 0;

    signal command_pos : integer range 1 to 6 := 1;
    signal byte_pos : integer range 1 to 17 := 1;

    signal state : integer range 1 to 22 := 1;


begin

    process(clk)
    begin
        if rising_edge(clk) then
            en_timing <= en_timing + 1;
            if en_timing <= 50000 then
                lcd_e <= '1';

            elsif (en_timing > 50000 and en_timing < 100000) then 
                lcd_e <= '0';

            elsif (en_timing = 100000) then
                en_timing <= 0;
				state <= state + 1;

                if(state <= 5) then
                    command_pos <= command_pos + 1;
                    
                elsif (state > 5) then
                    byte_pos <= byte_pos + 1;
                end if;
                
                if (state = 21) then
                    command_pos <= 5;
                    byte_pos <= 1;
                    state <= 5;
                end if;

            end if;


            if state <= 5 then      -- send command
                lcd_rw <= '0';
                lcd_rs <= '0';

                data_out <= command_rom(command_pos);


            elsif state > 5 then    -- send data
                lcd_rw <= '0';
                lcd_rs <= '1';

                data_out <= byte_in( (8*byte_pos)-1  downto  (8*byte_pos)-8 );

            end if;

        end if;

    end process;


end architecture arch;



 